----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    14:43:04 10/30/2016 
-- Design Name: 
-- Module Name:    PSR - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx primitives in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity PSR is
    Port ( ENTRADA_NZVC : in  STD_LOGIC_VECTOR (3 downto 0);
           RST : in  STD_LOGIC;
           CLK : in  STD_LOGIC;
           CARRY : out  STD_LOGIC;
			  ENTRADA_NCWP : in  STD_LOGIC;
			  SALIDA_CWP : out  STD_LOGIC);
end PSR;

architecture Behavioral of PSR is

begin
	process(ENTRADA_NZVC,RST,CLK,ENTRADA_NCWP)
	begin
		if RST='1' then
			SALIDA_CWP <= '0';
			CARRY <= '0';
		else
			if rising_edge(CLK) then
				if  ENTRADA_NCWP = '1' then
					 SALIDA_CWP <= '1';
				else
					SALIDA_CWP <= '0';
				end if;
				CARRY <= ENTRADA_NZVC(0);
			end if;
			
		end if;
	end process;

end Behavioral;

